module dayN

import util

pub fn solve_a(data string) !string {
    mut result := answer
    return result
}

pub fn solve_b(data string) !string {
    mut result := "answer"

    return result
}